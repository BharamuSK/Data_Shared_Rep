import uvm_pkg::*;      //uvm libraray files 
`include "uvm_macros.svh"//uvm librarty files `  they run during compilation time

`include "apb_tb.sv";
